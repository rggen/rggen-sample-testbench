class env_ral_model extends block_0_block_model #(
  .REGISTER_9           (block_1_block_model  ),
  .INTEGRATE_REGISTER_9 (1                    )
);
  `tue_object_default_constructor(env_ral_model)
  `uvm_object_utils(env_ral_model)
endclass
